library ieee;
use ieee.std_logic_1164.all;

entity sample_mem is 
	port (
		
	);